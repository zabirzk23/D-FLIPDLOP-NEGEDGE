module DFLIPFLOPNEGEDGE(D,Clock,Q,Qbar);
input D,Clock;
output reg Q,Qbar;
always @ // use negative edge clock for triggereing condition 
//compute D flipflop logic here
 endmodule
