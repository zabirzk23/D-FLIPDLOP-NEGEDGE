library verilog;
use verilog.vl_types.all;
entity DFLIPFLOPNEGEDGE_vlg_vec_tst is
end DFLIPFLOPNEGEDGE_vlg_vec_tst;
